module SumaPF_TB();

	//signals
	logic [31:0] a;
	logic [31:0] b;
	logic [31:0] result;
			  
	//DUT instance
	SumaPF DUT(a,b,result);
	
	//Test
	initial begin	
	a = 32'b11000010110010001000000000000000;//-100.25
	b = 32'b11000011100110001100100010110100;//-305.568
	#10;
	a = 32'b01000001101000100110011001100110;//20.3
	b = 32'b01000100000011100100000110101010;//50.263
	#10;
	a = 32'b01000010111100000000101000111101;//120.02
	b = 32'b01000100011110100001011110001101;//1000.368
	#10;
	a = 32'b11000010111100000000101000111101;//-120.02
	b = 32'b11000100000011100100000110101010;//-569.026
	#10;
	a = 32'b01000011010010001110010011000011;//200.8936
	b = 32'b01000011010010010100001010101010;//201.2604
	#10;
	a = 32'b01000010111100000000101000111101;//120.02
	b = 32'b01000100000011100100000110101010;//569.026
	#10;
	a = 32'b11000100011110100001011110001101;//-1000.368
	b = 32'b11000100000011100100000110101010;//-50.263
	#10;
	a = 32'b01000010111100000000101000111101;//120.02
	b = 32'b01000100000011100100000110101010;//569.026
	#10;
	 
	end

endmodule
