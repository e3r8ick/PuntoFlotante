module sumaPF